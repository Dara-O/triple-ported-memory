`ifndef _SHARED_PARAMS_
`define _SHARED_PARAMS_
// PARAMETERS FOR THE DIFFERENT PORT PRIORITIES
parameter PRIORITY_123 = 0;
parameter PRIORITY_132 = 1;
parameter PRIORITY_213 = 2;
parameter PRIORITY_231 = 3;
parameter PRIORITY_312 = 4;
parameter PRIORITY_321 = 5;

// PARAMETERS FOR IDENTIFYING THE ORIGINAL PORT OF A REORDERED PRIORITY PORT
parameter ORIG_PORT_1_ID = 1;
parameter ORIG_PORT_2_ID = 2;
parameter ORIG_PORT_3_ID = 3;
`endif